//this module is a tree based comparator